module Equiv_RecF32ToF32(
    input [32:0] io_in,
    output[31:0] io_out,
    output io_isBadNaN,
    output[8:0] io_smallExp,
    output io_goodExp
);

  wire T0;
  wire T1;
  wire[22:0] T2;
  wire T3;
  wire T4;
  wire[8:0] smallExp;
  wire[32:0] T5;
  wire[28:0] T6;
  wire[22:0] T7;
  wire[24:0] T8;
  wire[24:0] T9;
  wire[23:0] T10;
  wire[22:0] T11;
  wire[21:0] T12;
  wire[44:0] T13;
  wire[5:0] T15;
  wire[9:0] T16;
  wire[9:0] T17;
  wire[9:0] T18;
  wire[8:0] T19;
  wire[8:0] T20;
  wire[8:0] T21;
  wire[8:0] T76;
  wire[3:0] T22;
  wire[2:0] T23;
  wire[2:0] T77;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire[2:0] T27;
  wire[2:0] T28;
  wire T29;
  wire T30;
  wire[8:0] T31;
  wire T32;
  wire T33;
  wire[23:0] T34;
  wire T35;
  wire[2:0] T36;
  wire[31:0] T37;
  wire[30:0] T38;
  wire[22:0] T39;
  wire[22:0] T40;
  wire[22:0] T41;
  wire[24:0] T42;
  wire[24:0] T43;
  wire[23:0] T44;
  wire[22:0] T45;
  wire T46;
  wire T47;
  wire[2:0] T48;
  wire[8:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[1:0] T55;
  wire[22:0] T56;
  wire[23:0] T57;
  wire[4:0] T58;
  wire[4:0] T59;
  wire[9:0] T60;
  wire[9:0] T61;
  wire[9:0] T62;
  wire[23:0] T63;
  wire T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T78;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire[7:0] T73;
  wire T74;
  wire T75;


  assign io_goodExp = T0;
  assign T0 = T3 | T1;
  assign T1 = T2 == 23'h0;
  assign T2 = io_in[22:0];
  assign T3 = T4 ^ 1'h1;
  assign T4 = T31 < smallExp;
  assign smallExp = T5[31:23];
  assign T5 = {T22, T6};
  assign T6 = {T15, T7};
  assign T7 = T8[22:0];
  assign T8 = T9;
  assign T9 = {1'h0, T10};
  assign T10 = {1'h1, T11};
  assign T11 = T12 << 1'h1;
  assign T12 = T13[21:0];
  assign T13 = 23'h1 << 5'h16;
  assign T15 = T16[5:0];
  assign T16 = T17;
  assign T17 = T18;
  assign T18 = {1'h0, T19};
  assign T19 = T20;
  assign T20 = T21 + 9'h82;
  assign T21 = T76 ^ 9'h1ff;
  assign T76 = {4'h0, 5'h16};
  assign T22 = {T30, T23};
  assign T23 = T27 | T77;
  assign T77 = {2'h0, T24};
  assign T24 = T25;
  assign T25 = T26 == 2'h3;
  assign T26 = T20[8:7];
  assign T27 = T29 ? 3'h0 : T28;
  assign T28 = T16[8:6];
  assign T29 = 1'h0;
  assign T30 = 1'h0;
  assign T31 = io_in[31:23];
  assign io_smallExp = smallExp;
  assign io_isBadNaN = T32;
  assign T32 = T35 & T33;
  assign T33 = T34 != 24'hffffff;
  assign T34 = io_in[23:0];
  assign T35 = T36 == 3'h7;
  assign T36 = io_in[31:29];
  assign io_out = T37;
  assign T37 = {T74, T38};
  assign T38 = {T65, T39};
  assign T39 = T64 ? T56 : T40;
  assign T40 = T50 ? 23'h0 : T41;
  assign T41 = T42[22:0];
  assign T42 = T43;
  assign T43 = {1'h0, T44};
  assign T44 = {T46, T45};
  assign T45 = io_in[22:0];
  assign T46 = T47 ^ 1'h1;
  assign T47 = T48 == 3'h0;
  assign T48 = T49[8:6];
  assign T49 = io_in[31:23];
  assign T50 = T51;
  assign T51 = T54 & T52;
  assign T52 = T53 ^ 1'h1;
  assign T53 = T49[6];
  assign T54 = T55 == 2'h3;
  assign T55 = T49[8:7];
  assign T56 = T57[22:0];
  assign T57 = T63 >> T58;
  assign T58 = 5'h1 - T59;
  assign T59 = T60[4:0];
  assign T60 = T61;
  assign T61 = T62;
  assign T62 = {1'h0, T49};
  assign T63 = T42 >> 1'h1;
  assign T64 = $signed(T60) < $signed(9'h82);
  assign T65 = T71 | T66;
  assign T66 = 8'h0 - T78;
  assign T78 = {7'h0, T67};
  assign T67 = T68 | T50;
  assign T68 = T69;
  assign T69 = T54 & T70;
  assign T70 = T49[6];
  assign T71 = T64 ? 8'h0 : T72;
  assign T72 = T73 - 8'h81;
  assign T73 = T60[7:0];
  assign T74 = T75;
  assign T75 = io_in[32];
endmodule

