module Equiv_RecF32ToF32(
    input [32:0] io_in,
    output[31:0] io_out,
    output io_isZeroGood,
    output io_isBadExp,
    output io_isSubnormalGood
);

  wire T0;
  wire T1;
  wire[8:0] numZeros;
  wire[8:0] exp;
  wire[8:0] T140;
  wire[4:0] T141;
  wire[4:0] T142;
  wire[4:0] T143;
  wire[4:0] T144;
  wire[4:0] T145;
  wire[4:0] T146;
  wire[4:0] T147;
  wire[4:0] T148;
  wire[4:0] T149;
  wire[4:0] T150;
  wire[4:0] T151;
  wire[4:0] T152;
  wire[4:0] T153;
  wire[4:0] T154;
  wire[4:0] T155;
  wire[4:0] T156;
  wire[4:0] T157;
  wire[4:0] T158;
  wire[4:0] T159;
  wire[4:0] T160;
  wire[4:0] T161;
  wire[4:0] T162;
  wire T163;
  wire[22:0] T3;
  wire[6:0] T4;
  wire[2:0] T5;
  wire T6;
  wire[2:0] T7;
  wire[6:0] T8;
  wire[22:0] T9;
  wire[6:0] T10;
  wire[2:0] T11;
  wire T12;
  wire[2:0] T13;
  wire[6:0] T14;
  wire[22:0] sig;
  wire[1:0] T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire[3:0] T19;
  wire[1:0] T20;
  wire T21;
  wire[1:0] T22;
  wire[3:0] T23;
  wire T24;
  wire[1:0] T25;
  wire T26;
  wire[1:0] T27;
  wire T28;
  wire[15:0] T29;
  wire[15:0] T30;
  wire[15:0] T31;
  wire[14:0] T32;
  wire[15:0] T33;
  wire[15:0] T34;
  wire[15:0] T35;
  wire[13:0] T36;
  wire[15:0] T37;
  wire[15:0] T38;
  wire[15:0] T39;
  wire[11:0] T40;
  wire[15:0] T41;
  wire[15:0] T42;
  wire[15:0] T43;
  wire[7:0] T44;
  wire[15:0] T45;
  wire[15:0] T46;
  wire[15:0] T164;
  wire[7:0] T47;
  wire[15:0] T48;
  wire[15:0] T165;
  wire[11:0] T49;
  wire[15:0] T50;
  wire[15:0] T166;
  wire[13:0] T51;
  wire[15:0] T52;
  wire[15:0] T167;
  wire[14:0] T53;
  wire[1:0] T54;
  wire T55;
  wire[1:0] T56;
  wire T57;
  wire[3:0] T58;
  wire[1:0] T59;
  wire T60;
  wire[1:0] T61;
  wire[3:0] T62;
  wire T63;
  wire[1:0] T64;
  wire T65;
  wire[1:0] T66;
  wire T67;
  wire[15:0] T68;
  wire[15:0] T69;
  wire[15:0] T70;
  wire[14:0] T71;
  wire[15:0] T72;
  wire[15:0] T73;
  wire[15:0] T74;
  wire[13:0] T75;
  wire[15:0] T76;
  wire[15:0] T77;
  wire[15:0] T78;
  wire[11:0] T79;
  wire[15:0] T80;
  wire[15:0] T81;
  wire[15:0] T82;
  wire[7:0] T83;
  wire[15:0] T84;
  wire[15:0] T85;
  wire[15:0] T168;
  wire[7:0] T86;
  wire[15:0] T87;
  wire[15:0] T169;
  wire[11:0] T88;
  wire[15:0] T89;
  wire[15:0] T170;
  wire[13:0] T90;
  wire[15:0] T91;
  wire[15:0] T171;
  wire[14:0] T92;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire isSubnormal;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire[2:0] exp3;
  wire T98;
  wire T99;
  wire T100;
  wire[31:0] T101;
  wire[30:0] T102;
  wire[22:0] T103;
  wire[22:0] T104;
  wire[22:0] T105;
  wire[24:0] T106;
  wire[24:0] T107;
  wire[23:0] T108;
  wire[22:0] T109;
  wire T110;
  wire T111;
  wire[2:0] T112;
  wire[8:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire[1:0] T119;
  wire[22:0] T120;
  wire[23:0] T121;
  wire[4:0] T122;
  wire[4:0] T123;
  wire[9:0] T124;
  wire[9:0] T125;
  wire[9:0] T126;
  wire[23:0] T127;
  wire T128;
  wire[7:0] T129;
  wire[7:0] T130;
  wire[7:0] T193;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire[7:0] T135;
  wire[7:0] T136;
  wire[7:0] T137;
  wire T138;
  wire T139;


  assign io_isSubnormalGood = T0;
  assign T0 = isSubnormal & T1;
  assign T1 = T140 == numZeros;
  assign numZeros = exp - 9'h82;
  assign exp = io_in[31:23];
  assign T140 = {4'h0, T141};
  assign T141 = T192 ? 1'h0 : T142;
  assign T142 = T191 ? 1'h1 : T143;
  assign T143 = T190 ? 2'h2 : T144;
  assign T144 = T189 ? 2'h3 : T145;
  assign T145 = T188 ? 3'h4 : T146;
  assign T146 = T187 ? 3'h5 : T147;
  assign T147 = T186 ? 3'h6 : T148;
  assign T148 = T185 ? 3'h7 : T149;
  assign T149 = T184 ? 4'h8 : T150;
  assign T150 = T183 ? 4'h9 : T151;
  assign T151 = T182 ? 4'ha : T152;
  assign T152 = T181 ? 4'hb : T153;
  assign T153 = T180 ? 4'hc : T154;
  assign T154 = T179 ? 4'hd : T155;
  assign T155 = T178 ? 4'he : T156;
  assign T156 = T177 ? 4'hf : T157;
  assign T157 = T176 ? 5'h10 : T158;
  assign T158 = T175 ? 5'h11 : T159;
  assign T159 = T174 ? 5'h12 : T160;
  assign T160 = T173 ? 5'h13 : T161;
  assign T161 = T172 ? 5'h14 : T162;
  assign T162 = T163 ? 5'h15 : 5'h16;
  assign T163 = T3[21];
  assign T3 = {T68, T4};
  assign T4 = {T58, T5};
  assign T5 = {T54, T6};
  assign T6 = T7[2];
  assign T7 = T8[6:4];
  assign T8 = T9[22:16];
  assign T9 = {T29, T10};
  assign T10 = {T19, T11};
  assign T11 = {T15, T12};
  assign T12 = T13[2];
  assign T13 = T14[6:4];
  assign T14 = sig[22:16];
  assign sig = io_in[22:0];
  assign T15 = {T18, T16};
  assign T16 = T17[1];
  assign T17 = T13[1:0];
  assign T18 = T17[0];
  assign T19 = {T25, T20};
  assign T20 = {T24, T21};
  assign T21 = T22[1];
  assign T22 = T23[3:2];
  assign T23 = T14[3:0];
  assign T24 = T22[0];
  assign T25 = {T28, T26};
  assign T26 = T27[1];
  assign T27 = T23[1:0];
  assign T28 = T27[0];
  assign T29 = T52 | T30;
  assign T30 = T31 & 16'haaaa;
  assign T31 = T32 << 1'h1;
  assign T32 = T33[14:0];
  assign T33 = T50 | T34;
  assign T34 = T35 & 16'hcccc;
  assign T35 = T36 << 2'h2;
  assign T36 = T37[13:0];
  assign T37 = T48 | T38;
  assign T38 = T39 & 16'hf0f0;
  assign T39 = T40 << 3'h4;
  assign T40 = T41[11:0];
  assign T41 = T46 | T42;
  assign T42 = T43 & 16'hff00;
  assign T43 = T44 << 4'h8;
  assign T44 = T45[7:0];
  assign T45 = sig[15:0];
  assign T46 = T164 & 16'hff;
  assign T164 = {8'h0, T47};
  assign T47 = T45 >> 4'h8;
  assign T48 = T165 & 16'hf0f;
  assign T165 = {4'h0, T49};
  assign T49 = T41 >> 3'h4;
  assign T50 = T166 & 16'h3333;
  assign T166 = {2'h0, T51};
  assign T51 = T37 >> 2'h2;
  assign T52 = T167 & 16'h5555;
  assign T167 = {1'h0, T53};
  assign T53 = T33 >> 1'h1;
  assign T54 = {T57, T55};
  assign T55 = T56[1];
  assign T56 = T7[1:0];
  assign T57 = T56[0];
  assign T58 = {T64, T59};
  assign T59 = {T63, T60};
  assign T60 = T61[1];
  assign T61 = T62[3:2];
  assign T62 = T8[3:0];
  assign T63 = T61[0];
  assign T64 = {T67, T65};
  assign T65 = T66[1];
  assign T66 = T62[1:0];
  assign T67 = T66[0];
  assign T68 = T91 | T69;
  assign T69 = T70 & 16'haaaa;
  assign T70 = T71 << 1'h1;
  assign T71 = T72[14:0];
  assign T72 = T89 | T73;
  assign T73 = T74 & 16'hcccc;
  assign T74 = T75 << 2'h2;
  assign T75 = T76[13:0];
  assign T76 = T87 | T77;
  assign T77 = T78 & 16'hf0f0;
  assign T78 = T79 << 3'h4;
  assign T79 = T80[11:0];
  assign T80 = T85 | T81;
  assign T81 = T82 & 16'hff00;
  assign T82 = T83 << 4'h8;
  assign T83 = T84[7:0];
  assign T84 = T9[15:0];
  assign T85 = T168 & 16'hff;
  assign T168 = {8'h0, T86};
  assign T86 = T84 >> 4'h8;
  assign T87 = T169 & 16'hf0f;
  assign T169 = {4'h0, T88};
  assign T88 = T80 >> 3'h4;
  assign T89 = T170 & 16'h3333;
  assign T170 = {2'h0, T90};
  assign T90 = T76 >> 2'h2;
  assign T91 = T171 & 16'h5555;
  assign T171 = {1'h0, T92};
  assign T92 = T72 >> 1'h1;
  assign T172 = T3[20];
  assign T173 = T3[19];
  assign T174 = T3[18];
  assign T175 = T3[17];
  assign T176 = T3[16];
  assign T177 = T3[15];
  assign T178 = T3[14];
  assign T179 = T3[13];
  assign T180 = T3[12];
  assign T181 = T3[11];
  assign T182 = T3[10];
  assign T183 = T3[9];
  assign T184 = T3[8];
  assign T185 = T3[7];
  assign T186 = T3[6];
  assign T187 = T3[5];
  assign T188 = T3[4];
  assign T189 = T3[3];
  assign T190 = T3[2];
  assign T191 = T3[1];
  assign T192 = T3[0];
  assign isSubnormal = T94 & T93;
  assign T93 = 9'h6b <= exp;
  assign T94 = exp < 9'h82;
  assign io_isBadExp = T95;
  assign T95 = T97 & T96;
  assign T96 = exp < 9'h6b;
  assign T97 = exp3 != 3'h0;
  assign exp3 = exp[8:6];
  assign io_isZeroGood = T98;
  assign T98 = T100 | T99;
  assign T99 = sig == 23'h0;
  assign T100 = exp3 != 3'h0;
  assign io_out = T101;
  assign T101 = {T138, T102};
  assign T102 = {T129, T103};
  assign T103 = T128 ? T120 : T104;
  assign T104 = T114 ? 23'h0 : T105;
  assign T105 = T106[22:0];
  assign T106 = T107;
  assign T107 = {1'h0, T108};
  assign T108 = {T110, T109};
  assign T109 = io_in[22:0];
  assign T110 = T111 ^ 1'h1;
  assign T111 = T112 == 3'h0;
  assign T112 = T113[8:6];
  assign T113 = io_in[31:23];
  assign T114 = T115;
  assign T115 = T118 & T116;
  assign T116 = T117 ^ 1'h1;
  assign T117 = T113[6];
  assign T118 = T119 == 2'h3;
  assign T119 = T113[8:7];
  assign T120 = T121[22:0];
  assign T121 = T127 >> T122;
  assign T122 = 5'h1 - T123;
  assign T123 = T124[4:0];
  assign T124 = T125;
  assign T125 = T126;
  assign T126 = {1'h0, T113};
  assign T127 = T106 >> 1'h1;
  assign T128 = $signed(T124) < $signed(9'h82);
  assign T129 = T135 | T130;
  assign T130 = 8'h0 - T193;
  assign T193 = {7'h0, T131};
  assign T131 = T132 | T114;
  assign T132 = T133;
  assign T133 = T118 & T134;
  assign T134 = T113[6];
  assign T135 = T128 ? 8'h0 : T136;
  assign T136 = T137 - 8'h81;
  assign T137 = T124[7:0];
  assign T138 = T139;
  assign T139 = io_in[32];
endmodule

